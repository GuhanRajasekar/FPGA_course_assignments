`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12.04.2024 19:48:13
// Design Name: 
// Module Name: cordic_tanh_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cordic_tanh_tb;
reg clk, rst;
reg signed  [19:0] target_angle;
wire signed [19:0] tanh;

cordic_tanh balout(.clk(clk), .rst(rst), .target_angle(target_angle), .tanh(tanh));

always #2 clk = ~clk;
initial
  begin
    #0 clk = 1'b1; rst = 1'b0;
    #2 rst = 1'b1;

#15 target_angle = 20'b11111110110000000000; //-5.0 radians
#15 target_angle = 20'b11111110110000110100; //-4.949748743718593 radians
#15 target_angle = 20'b11111110110001100111; //-4.899497487437186 radians
#15 target_angle = 20'b11111110110010011011; //-4.849246231155779 radians
#15 target_angle = 20'b11111110110011001110; //-4.798994974874372 radians
#15 target_angle = 20'b11111110110100000010; //-4.748743718592965 radians
#15 target_angle = 20'b11111110110100110101; //-4.698492462311558 radians
#15 target_angle = 20'b11111110110101101001; //-4.648241206030151 radians
#15 target_angle = 20'b11111110110110011100; //-4.597989949748744 radians
#15 target_angle = 20'b11111110110111010000; //-4.547738693467337 radians
#15 target_angle = 20'b11111110111000000011; //-4.49748743718593 radians
#15 target_angle = 20'b11111110111000110111; //-4.447236180904523 radians
#15 target_angle = 20'b11111110111001101010; //-4.396984924623116 radians
#15 target_angle = 20'b11111110111010011101; //-4.346733668341709 radians
#15 target_angle = 20'b11111110111011010001; //-4.296482412060302 radians
#15 target_angle = 20'b11111110111100000100; //-4.2462311557788945 radians
#15 target_angle = 20'b11111110111100111000; //-4.1959798994974875 radians
#15 target_angle = 20'b11111110111101101011; //-4.1457286432160805 radians
#15 target_angle = 20'b11111110111110011111; //-4.0954773869346734 radians
#15 target_angle = 20'b11111110111111010010; //-4.045226130653266 radians
#15 target_angle = 20'b11111111000000000110; //-3.9949748743718594 radians
#15 target_angle = 20'b11111111000000111001; //-3.9447236180904524 radians
#15 target_angle = 20'b11111111000001101101; //-3.8944723618090453 radians
#15 target_angle = 20'b11111111000010100000; //-3.8442211055276383 radians
#15 target_angle = 20'b11111111000011010011; //-3.7939698492462313 radians
#15 target_angle = 20'b11111111000100000111; //-3.7437185929648242 radians
#15 target_angle = 20'b11111111000100111010; //-3.693467336683417 radians
#15 target_angle = 20'b11111111000101101110; //-3.64321608040201 radians
#15 target_angle = 20'b11111111000110100001; //-3.592964824120603 radians
#15 target_angle = 20'b11111111000111010101; //-3.542713567839196 radians
#15 target_angle = 20'b11111111001000001000; //-3.492462311557789 radians
#15 target_angle = 20'b11111111001000111100; //-3.442211055276382 radians
#15 target_angle = 20'b11111111001001101111; //-3.391959798994975 radians
#15 target_angle = 20'b11111111001010100011; //-3.341708542713568 radians
#15 target_angle = 20'b11111111001011010110; //-3.291457286432161 radians
#15 target_angle = 20'b11111111001100001010; //-3.241206030150754 radians
#15 target_angle = 20'b11111111001100111101; //-3.190954773869347 radians
#15 target_angle = 20'b11111111001101110000; //-3.14070351758794 radians
#15 target_angle = 20'b11111111001110100100; //-3.090452261306533 radians
#15 target_angle = 20'b11111111001111010111; //-3.040201005025126 radians
#15 target_angle = 20'b11111111010000001011; //-2.9899497487437183 radians
#15 target_angle = 20'b11111111010000111110; //-2.9396984924623113 radians
#15 target_angle = 20'b11111111010001110010; //-2.8894472361809043 radians
#15 target_angle = 20'b11111111010010100101; //-2.8391959798994972 radians
#15 target_angle = 20'b11111111010011011001; //-2.78894472361809 radians
#15 target_angle = 20'b11111111010100001100; //-2.738693467336683 radians
#15 target_angle = 20'b11111111010101000000; //-2.688442211055276 radians
#15 target_angle = 20'b11111111010101110011; //-2.638190954773869 radians
#15 target_angle = 20'b11111111010110100110; //-2.587939698492462 radians
#15 target_angle = 20'b11111111010111011010; //-2.537688442211055 radians
#15 target_angle = 20'b11111111011000001101; //-2.487437185929648 radians
#15 target_angle = 20'b11111111011001000001; //-2.437185929648241 radians
#15 target_angle = 20'b11111111011001110100; //-2.386934673366834 radians
#15 target_angle = 20'b11111111011010101000; //-2.336683417085427 radians
#15 target_angle = 20'b11111111011011011011; //-2.28643216080402 radians
#15 target_angle = 20'b11111111011100001111; //-2.236180904522613 radians
#15 target_angle = 20'b11111111011101000010; //-2.185929648241206 radians
#15 target_angle = 20'b11111111011101110110; //-2.135678391959799 radians
#15 target_angle = 20'b11111111011110101001; //-2.0854271356783918 radians
#15 target_angle = 20'b11111111011111011100; //-2.0351758793969847 radians
#15 target_angle = 20'b11111111100000010000; //-1.9849246231155777 radians
#15 target_angle = 20'b11111111100001000011; //-1.9346733668341707 radians
#15 target_angle = 20'b11111111100001110111; //-1.8844221105527637 radians
#15 target_angle = 20'b11111111100010101010; //-1.8341708542713566 radians
#15 target_angle = 20'b11111111100011011110; //-1.7839195979899496 radians
#15 target_angle = 20'b11111111100100010001; //-1.7336683417085426 radians
#15 target_angle = 20'b11111111100101000101; //-1.6834170854271355 radians
#15 target_angle = 20'b11111111100101111000; //-1.6331658291457285 radians
#15 target_angle = 20'b11111111100110101100; //-1.5829145728643215 radians
#15 target_angle = 20'b11111111100111011111; //-1.5326633165829144 radians
#15 target_angle = 20'b11111111101000010011; //-1.4824120603015074 radians
#15 target_angle = 20'b11111111101001000110; //-1.4321608040201004 radians
#15 target_angle = 20'b11111111101001111001; //-1.3819095477386933 radians
#15 target_angle = 20'b11111111101010101101; //-1.3316582914572863 radians
#15 target_angle = 20'b11111111101011100000; //-1.2814070351758793 radians
#15 target_angle = 20'b11111111101100010100; //-1.2311557788944723 radians
#15 target_angle = 20'b11111111101101000111; //-1.1809045226130652 radians
#15 target_angle = 20'b11111111101101111011; //-1.1306532663316582 radians
#15 target_angle = 20'b11111111101110101110; //-1.0804020100502512 radians
#15 target_angle = 20'b11111111101111100010; //-1.0301507537688441 radians
#15 target_angle = 20'b11111111110000010101; //-0.9798994974874367 radians
#15 target_angle = 20'b11111111110001001001; //-0.9296482412060296 radians
#15 target_angle = 20'b11111111110001111100; //-0.8793969849246226 radians
#15 target_angle = 20'b11111111110010101111; //-0.8291457286432156 radians
#15 target_angle = 20'b11111111110011100011; //-0.7788944723618085 radians
#15 target_angle = 20'b11111111110100010110; //-0.7286432160804015 radians
#15 target_angle = 20'b11111111110101001010; //-0.6783919597989945 radians
#15 target_angle = 20'b11111111110101111101; //-0.6281407035175874 radians
#15 target_angle = 20'b11111111110110110001; //-0.5778894472361804 radians
#15 target_angle = 20'b11111111110111100100; //-0.5276381909547734 radians
#15 target_angle = 20'b11111111111000011000; //-0.47738693467336635 radians
#15 target_angle = 20'b11111111111001001011; //-0.4271356783919593 radians
#15 target_angle = 20'b11111111111001111111; //-0.3768844221105523 radians
#15 target_angle = 20'b11111111111010110010; //-0.32663316582914526 radians
#15 target_angle = 20'b11111111111011100101; //-0.2763819095477382 radians
#15 target_angle = 20'b11111111111100011001; //-0.2261306532663312 radians
#15 target_angle = 20'b11111111111101001100; //-0.17587939698492416 radians
#15 target_angle = 20'b11111111111110000000; //-0.12562814070351713 radians
#15 target_angle = 20'b11111111111110110011; //-0.0753768844221101 radians
#15 target_angle = 20'b11111111111111100111; //-0.02512562814070307 radians
#15 target_angle = 20'b00000000000000011001; //0.02512562814070396 radians
#15 target_angle = 20'b00000000000001001101; //0.07537688442211099 radians
#15 target_angle = 20'b00000000000010000000; //0.12562814070351802 radians
#15 target_angle = 20'b00000000000010110100; //0.17587939698492505 radians
#15 target_angle = 20'b00000000000011100111; //0.22613065326633208 radians
#15 target_angle = 20'b00000000000100011011; //0.2763819095477391 radians
#15 target_angle = 20'b00000000000101001110; //0.32663316582914614 radians
#15 target_angle = 20'b00000000000110000001; //0.3768844221105532 radians
#15 target_angle = 20'b00000000000110110101; //0.4271356783919602 radians
#15 target_angle = 20'b00000000000111101000; //0.47738693467336724 radians
#15 target_angle = 20'b00000000001000011100; //0.5276381909547743 radians
#15 target_angle = 20'b00000000001001001111; //0.5778894472361813 radians
#15 target_angle = 20'b00000000001010000011; //0.6281407035175883 radians
#15 target_angle = 20'b00000000001010110110; //0.6783919597989954 radians
#15 target_angle = 20'b00000000001011101010; //0.7286432160804024 radians
#15 target_angle = 20'b00000000001100011101; //0.7788944723618094 radians
#15 target_angle = 20'b00000000001101010001; //0.8291457286432165 radians
#15 target_angle = 20'b00000000001110000100; //0.8793969849246235 radians
#15 target_angle = 20'b00000000001110110111; //0.9296482412060305 radians
#15 target_angle = 20'b00000000001111101011; //0.9798994974874375 radians
#15 target_angle = 20'b00000000010000011110; //1.0301507537688446 radians
#15 target_angle = 20'b00000000010001010010; //1.0804020100502516 radians
#15 target_angle = 20'b00000000010010000101; //1.1306532663316586 radians
#15 target_angle = 20'b00000000010010111001; //1.1809045226130657 radians
#15 target_angle = 20'b00000000010011101100; //1.2311557788944727 radians
#15 target_angle = 20'b00000000010100100000; //1.2814070351758797 radians
#15 target_angle = 20'b00000000010101010011; //1.3316582914572868 radians
#15 target_angle = 20'b00000000010110000111; //1.3819095477386938 radians
#15 target_angle = 20'b00000000010110111010; //1.4321608040201008 radians
#15 target_angle = 20'b00000000010111101101; //1.4824120603015079 radians
#15 target_angle = 20'b00000000011000100001; //1.5326633165829149 radians
#15 target_angle = 20'b00000000011001010100; //1.582914572864322 radians
#15 target_angle = 20'b00000000011010001000; //1.633165829145729 radians
#15 target_angle = 20'b00000000011010111011; //1.683417085427136 radians
#15 target_angle = 20'b00000000011011101111; //1.733668341708543 radians
#15 target_angle = 20'b00000000011100100010; //1.78391959798995 radians
#15 target_angle = 20'b00000000011101010110; //1.834170854271357 radians
#15 target_angle = 20'b00000000011110001001; //1.884422110552764 radians
#15 target_angle = 20'b00000000011110111101; //1.9346733668341711 radians
#15 target_angle = 20'b00000000011111110000; //1.9849246231155782 radians
#15 target_angle = 20'b00000000100000100100; //2.035175879396985 radians
#15 target_angle = 20'b00000000100001010111; //2.085427135678392 radians
#15 target_angle = 20'b00000000100010001010; //2.1356783919597992 radians
#15 target_angle = 20'b00000000100010111110; //2.1859296482412063 radians
#15 target_angle = 20'b00000000100011110001; //2.2361809045226133 radians
#15 target_angle = 20'b00000000100100100101; //2.2864321608040203 radians
#15 target_angle = 20'b00000000100101011000; //2.3366834170854274 radians
#15 target_angle = 20'b00000000100110001100; //2.3869346733668344 radians
#15 target_angle = 20'b00000000100110111111; //2.4371859296482414 radians
#15 target_angle = 20'b00000000100111110011; //2.4874371859296485 radians
#15 target_angle = 20'b00000000101000100110; //2.5376884422110555 radians
#15 target_angle = 20'b00000000101001011010; //2.5879396984924625 radians
#15 target_angle = 20'b00000000101010001101; //2.6381909547738696 radians
#15 target_angle = 20'b00000000101011000000; //2.6884422110552766 radians
#15 target_angle = 20'b00000000101011110100; //2.7386934673366836 radians
#15 target_angle = 20'b00000000101100100111; //2.7889447236180906 radians
#15 target_angle = 20'b00000000101101011011; //2.8391959798994977 radians
#15 target_angle = 20'b00000000101110001110; //2.8894472361809047 radians
#15 target_angle = 20'b00000000101111000010; //2.9396984924623117 radians
#15 target_angle = 20'b00000000101111110101; //2.9899497487437188 radians
#15 target_angle = 20'b00000000110000101001; //3.0402010050251267 radians
#15 target_angle = 20'b00000000110001011100; //3.090452261306533 radians
#15 target_angle = 20'b00000000110010010000; //3.1407035175879408 radians
#15 target_angle = 20'b00000000110011000011; //3.190954773869347 radians
#15 target_angle = 20'b00000000110011110110; //3.241206030150755 radians
#15 target_angle = 20'b00000000110100101010; //3.291457286432161 radians
#15 target_angle = 20'b00000000110101011101; //3.341708542713569 radians
#15 target_angle = 20'b00000000110110010001; //3.391959798994975 radians
#15 target_angle = 20'b00000000110111000100; //3.442211055276383 radians
#15 target_angle = 20'b00000000110111111000; //3.492462311557789 radians
#15 target_angle = 20'b00000000111000101011; //3.542713567839197 radians
#15 target_angle = 20'b00000000111001011111; //3.592964824120603 radians
#15 target_angle = 20'b00000000111010010010; //3.643216080402011 radians
#15 target_angle = 20'b00000000111011000110; //3.693467336683417 radians
#15 target_angle = 20'b00000000111011111001; //3.743718592964825 radians
#15 target_angle = 20'b00000000111100101101; //3.7939698492462313 radians
#15 target_angle = 20'b00000000111101100000; //3.844221105527639 radians
#15 target_angle = 20'b00000000111110010011; //3.8944723618090453 radians
#15 target_angle = 20'b00000000111111000111; //3.9447236180904532 radians
#15 target_angle = 20'b00000000111111111010; //3.9949748743718594 radians
#15 target_angle = 20'b00000001000000101110; //4.045226130653267 radians
#15 target_angle = 20'b00000001000001100001; //4.0954773869346734 radians
#15 target_angle = 20'b00000001000010010101; //4.145728643216081 radians
#15 target_angle = 20'b00000001000011001000; //4.1959798994974875 radians
#15 target_angle = 20'b00000001000011111100; //4.246231155778895 radians
#15 target_angle = 20'b00000001000100101111; //4.296482412060302 radians
#15 target_angle = 20'b00000001000101100011; //4.3467336683417095 radians
#15 target_angle = 20'b00000001000110010110; //4.396984924623116 radians
#15 target_angle = 20'b00000001000111001001; //4.4472361809045236 radians
#15 target_angle = 20'b00000001000111111101; //4.49748743718593 radians
#15 target_angle = 20'b00000001001000110000; //4.547738693467338 radians
#15 target_angle = 20'b00000001001001100100; //4.597989949748744 radians
#15 target_angle = 20'b00000001001010010111; //4.648241206030152 radians
#15 target_angle = 20'b00000001001011001011; //4.698492462311558 radians
#15 target_angle = 20'b00000001001011111110; //4.748743718592966 radians
#15 target_angle = 20'b00000001001100110010; //4.798994974874372 radians
#15 target_angle = 20'b00000001001101100101; //4.84924623115578 radians
#15 target_angle = 20'b00000001001110011001; //4.899497487437186 radians
#15 target_angle = 20'b00000001001111001100; //4.949748743718594 radians
#15 target_angle = 20'b00000001010000000000; //5.0 radians


      #50 $finish;
  end
endmodule
