`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 31.03.2024 12:50:29
// Design Name: 
// Module Name: cordic_tanh_inverse_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module cordic_tanh_inverse_tb;
  reg  signed  [19:0] y_input;
  reg  clk, rst;
  
  wire signed [19:0] z_res;
  
  cordic_tanh_inverse k(.clk(clk) , .rst(rst), .y_input(y_input), .z_res(z_res));
  
  always #2 clk = ~clk;
  
  initial 
     begin
      #0 clk = 1'b0; rst = 1'b0; 
      #1 rst = 1'b1;
//      #5 y_input = {{4'b1111},{16'b0000110011001101}} ; // y = -0.95
//      #5 y_input = {{4'b1111},{16'b0001100110011010}} ; // y = -0.9
//      #5 y_input = {{4'b1111},{16'b0010011001100111}} ; // y = -0.85
//      #5 y_input = {{4'b1111},{16'b0011001100110100}} ; // y = -0.8
//      #5 y_input = {{4'b1111},{16'b0100000000000000}} ; // y = -0.75
//      #5 y_input = {{4'b1111},{16'b0100110011001101}} ; // y = -0.7
//      #5 y_input = {{4'b1111},{16'b0101100110011010}} ; // y = -0.65
//      #5 y_input = {{4'b1111},{16'b0110011001100111}} ; // y = -0.6
//      #5 y_input = {{4'b1111},{16'b0111001100110100}} ; // y = -0.55
//      #5 y_input = {{4'b1111},{16'b1000000000000000}} ; // y = -0.5
//      #5 y_input = {{4'b1111},{16'b1000110011001101}} ; // y = -0.45
//      #5 y_input = {{4'b1111},{16'b1001100110011010}} ; // y = -0.4
//      #5 y_input = {{4'b1111},{16'b1010011001100111}} ; // y = -0.35
//      #5 y_input = {{4'b1111},{16'b1011001100110100}} ; // y = -0.3
//      #5 y_input = {{4'b1111},{16'b1100000000000000}} ; // y = -0.25
//      #5 y_input = {{4'b1111},{16'b1100110011001101}} ; // y = -0.2
//      #5 y_input = {{4'b1111},{16'b1101100110011010}} ; // y = -0.15
//      #5 y_input = {{4'b1111},{16'b1110011001100111}} ; // y = -0.1
//      #5 y_input = {{4'b1111},{16'b1111001100110100}} ; // y = -0.05
     
//      #5 y_input = {{4'b0000},{16'b0000000000000000}} ; // y = 0
//      #5 y_input = {{4'b0000},{16'b0000110011001100}} ; // y = 0.05
//      #5 y_input = {{4'b0000},{16'b0001100110011001}} ; // y = 0.1
//      #5 y_input = {{4'b0000},{16'b0010011001100110}} ; // y = 0.15
//      #5 y_input = {{4'b0000},{16'b0011001100110011}} ; // y = 0.2
//      #5 y_input = {{4'b0000},{16'b0100000000000000}} ; // y = 0.25
//      #5 y_input = {{4'b0000},{16'b0100110011001100}} ; // y = 0.3
//      #5 y_input = {{4'b0000},{16'b0101100110011001}} ; // y = 0.35
//      #5 y_input = {{4'b0000},{16'b0110011001100110}} ; // y = 0.4
//      #5 y_input = {{4'b0000},{16'b0111001100110011}} ; // y = 0.45
//      #5 y_input = {{4'b0000},{16'b1000000000000000}} ; // y = 0.5
//      #5 y_input = {{4'b0000},{16'b1000110011001100}} ; // y = 0.55
//      #5 y_input = {{4'b0000},{16'b1001100110011001}} ; // y = 0.6
//      #5 y_input = {{4'b0000},{16'b1010011001100110}} ; // y = 0.65
//      #5 y_input = {{4'b0000},{16'b1011001100110011}} ; // y = 0.7
//      #5 y_input = {{4'b0000},{16'b1100000000000000}} ; // y = 0.75
//      #5 y_input = {{4'b0000},{16'b1100110011001100}} ; // y = 0.8
//      #5 y_input = {{4'b0000},{16'b1101100110011001}} ; // y = 0.85
//      #5 y_input = {{4'b0000},{16'b1110011001100110}} ; // y = 0.9
//      #5 y_input = {{4'b0000},{16'b1111001100110011}} ; // y = 0.95
//      #5 y_input = {{4'b0001},{16'b0000000000000000}} ; // y = 0.95

#15 y_input = 20'b11110000110011001101; // y = -0.95 
#15 y_input = 20'b11110000111100111111; // y = -0.9404522613065326 
#15 y_input = 20'b11110001000110110001; // y = -0.9309045226130653 
#15 y_input = 20'b11110001010000100010; // y = -0.921356783919598 
#15 y_input = 20'b11110001011010010100; // y = -0.9118090452261306 
#15 y_input = 20'b11110001100100000110; // y = -0.9022613065326632 
#15 y_input = 20'b11110001101101111000; // y = -0.892713567839196 
#15 y_input = 20'b11110001110111101001; // y = -0.8831658291457286 
#15 y_input = 20'b11110010000001011011; // y = -0.8736180904522612 
#15 y_input = 20'b11110010001011001101; // y = -0.864070351758794 
#15 y_input = 20'b11110010010100111111; // y = -0.8545226130653266 
#15 y_input = 20'b11110010011110110000; // y = -0.8449748743718593 
#15 y_input = 20'b11110010101000100010; // y = -0.8354271356783919 
#15 y_input = 20'b11110010110010010100; // y = -0.8258793969849246 
#15 y_input = 20'b11110010111100000101; // y = -0.8163316582914573 
#15 y_input = 20'b11110011000101110111; // y = -0.8067839195979899 
#15 y_input = 20'b11110011001111101001; // y = -0.7972361809045225 
#15 y_input = 20'b11110011011001011011; // y = -0.7876884422110553 
#15 y_input = 20'b11110011100011001100; // y = -0.7781407035175879 
#15 y_input = 20'b11110011101100111110; // y = -0.7685929648241205 
#15 y_input = 20'b11110011110110110000; // y = -0.7590452261306533 
#15 y_input = 20'b11110100000000100001; // y = -0.7494974874371859 
#15 y_input = 20'b11110100001010010011; // y = -0.7399497487437185 
#15 y_input = 20'b11110100010100000101; // y = -0.7304020100502513 
#15 y_input = 20'b11110100011101110111; // y = -0.7208542713567839 
#15 y_input = 20'b11110100100111101000; // y = -0.7113065326633166 
#15 y_input = 20'b11110100110001011010; // y = -0.7017587939698492 
#15 y_input = 20'b11110100111011001100; // y = -0.6922110552763818 
#15 y_input = 20'b11110101000100111101; // y = -0.6826633165829146 
#15 y_input = 20'b11110101001110101111; // y = -0.6731155778894472 
#15 y_input = 20'b11110101011000100001; // y = -0.6635678391959798 
#15 y_input = 20'b11110101100010010011; // y = -0.6540201005025126 
#15 y_input = 20'b11110101101100000100; // y = -0.6444723618090452 
#15 y_input = 20'b11110101110101110110; // y = -0.6349246231155778 
#15 y_input = 20'b11110101111111101000; // y = -0.6253768844221106 
#15 y_input = 20'b11110110001001011010; // y = -0.6158291457286432 
#15 y_input = 20'b11110110010011001011; // y = -0.6062814070351759 
#15 y_input = 20'b11110110011100111101; // y = -0.5967336683417086 
#15 y_input = 20'b11110110100110101111; // y = -0.5871859296482411 
#15 y_input = 20'b11110110110000100000; // y = -0.5776381909547739 
#15 y_input = 20'b11110110111010010010; // y = -0.5680904522613065 
#15 y_input = 20'b11110111000100000100; // y = -0.5585427135678391 
#15 y_input = 20'b11110111001101110110; // y = -0.5489949748743719 
#15 y_input = 20'b11110111010111100111; // y = -0.5394472361809045 
#15 y_input = 20'b11110111100001011001; // y = -0.5298994974874371 
#15 y_input = 20'b11110111101011001011; // y = -0.5203517587939699 
#15 y_input = 20'b11110111110100111100; // y = -0.5108040201005025 
#15 y_input = 20'b11110111111110101110; // y = -0.5012562814070352 
#15 y_input = 20'b11111000001000100000; // y = -0.49170854271356784 
#15 y_input = 20'b11111000010010010010; // y = -0.48216080402010053 
#15 y_input = 20'b11111000011100000011; // y = -0.47261306532663316 
#15 y_input = 20'b11111000100101110101; // y = -0.46306532663316585 
#15 y_input = 20'b11111000101111100111; // y = -0.4535175879396985 
#15 y_input = 20'b11111000111001011000; // y = -0.4439698492462312 
#15 y_input = 20'b11111001000011001010; // y = -0.4344221105527638 
#15 y_input = 20'b11111001001100111100; // y = -0.42487437185929644 
#15 y_input = 20'b11111001010110101110; // y = -0.4153266331658292 
#15 y_input = 20'b11111001100000011111; // y = -0.4057788944723618 
#15 y_input = 20'b11111001101010010001; // y = -0.39623115577889445 
#15 y_input = 20'b11111001110100000011; // y = -0.3866834170854272 
#15 y_input = 20'b11111001111101110101; // y = -0.3771356783919598 
#15 y_input = 20'b11111010000111100110; // y = -0.36758793969849246 
#15 y_input = 20'b11111010010001011000; // y = -0.3580402010050251 
#15 y_input = 20'b11111010011011001010; // y = -0.34849246231155784 
#15 y_input = 20'b11111010100100111011; // y = -0.33894472361809047 
#15 y_input = 20'b11111010101110101101; // y = -0.3293969849246231 
#15 y_input = 20'b11111010111000011111; // y = -0.31984924623115585 
#15 y_input = 20'b11111011000010010001; // y = -0.3103015075376885 
#15 y_input = 20'b11111011001100000010; // y = -0.3007537688442211 
#15 y_input = 20'b11111011010101110100; // y = -0.29120603015075375 
#15 y_input = 20'b11111011011111100110; // y = -0.2816582914572865 
#15 y_input = 20'b11111011101001010111; // y = -0.2721105527638191 
#15 y_input = 20'b11111011110011001001; // y = -0.26256281407035176 
#15 y_input = 20'b11111011111100111011; // y = -0.2530150753768845 
#15 y_input = 20'b11111100000110101101; // y = -0.24346733668341713 
#15 y_input = 20'b11111100010000011110; // y = -0.23391959798994977 
#15 y_input = 20'b11111100011010010000; // y = -0.2243718592964824 
#15 y_input = 20'b11111100100100000010; // y = -0.21482412060301515 
#15 y_input = 20'b11111100101101110100; // y = -0.20527638190954778 
#15 y_input = 20'b11111100110111100101; // y = -0.1957286432160804 
#15 y_input = 20'b11111101000001010111; // y = -0.18618090452261304 
#15 y_input = 20'b11111101001011001001; // y = -0.1766331658291458 
#15 y_input = 20'b11111101010100111010; // y = -0.16708542713567842 
#15 y_input = 20'b11111101011110101100; // y = -0.15753768844221105 
#15 y_input = 20'b11111101101000011110; // y = -0.1479899497487438 
#15 y_input = 20'b11111101110010010000; // y = -0.13844221105527643 
#15 y_input = 20'b11111101111100000001; // y = -0.12889447236180906 
#15 y_input = 20'b11111110000101110011; // y = -0.1193467336683417 
#15 y_input = 20'b11111110001111100101; // y = -0.10979899497487444 
#15 y_input = 20'b11111110011001010110; // y = -0.10025125628140708 
#15 y_input = 20'b11111110100011001000; // y = -0.09070351758793971 
#15 y_input = 20'b11111110101100111010; // y = -0.08115577889447245 
#15 y_input = 20'b11111110110110101100; // y = -0.07160804020100509 
#15 y_input = 20'b11111111000000011101; // y = -0.06206030150753772 
#15 y_input = 20'b11111111001010001111; // y = -0.05251256281407035 
#15 y_input = 20'b11111111010100000001; // y = -0.042964824120603096 
#15 y_input = 20'b11111111011101110010; // y = -0.03341708542713573 
#15 y_input = 20'b11111111100111100100; // y = -0.023869346733668362 
#15 y_input = 20'b11111111110001010110; // y = -0.014321608040201106 
#15 y_input = 20'b11111111111011001000; // y = -0.004773869346733739 
#15 y_input = 20'b00000000000100111000; // y = 0.004773869346733628 
#15 y_input = 20'b00000000001110101010; // y = 0.014321608040200995 
#15 y_input = 20'b00000000011000011100; // y = 0.02386934673366825 
#15 y_input = 20'b00000000100010001110; // y = 0.03341708542713562 
#15 y_input = 20'b00000000101011111111; // y = 0.042964824120602985 
#15 y_input = 20'b00000000110101110001; // y = 0.05251256281407035 
#15 y_input = 20'b00000000111111100011; // y = 0.06206030150753761 
#15 y_input = 20'b00000001001001010100; // y = 0.07160804020100486 
#15 y_input = 20'b00000001010011000110; // y = 0.08115577889447234 
#15 y_input = 20'b00000001011100111000; // y = 0.0907035175879396 
#15 y_input = 20'b00000001100110101010; // y = 0.10025125628140708 
#15 y_input = 20'b00000001110000011011; // y = 0.10979899497487433 
#15 y_input = 20'b00000001111010001101; // y = 0.11934673366834159 
#15 y_input = 20'b00000010000011111111; // y = 0.12889447236180906 
#15 y_input = 20'b00000010001101110000; // y = 0.13844221105527632 
#15 y_input = 20'b00000010010111100010; // y = 0.14798994974874358 
#15 y_input = 20'b00000010100001010100; // y = 0.15753768844221105 
#15 y_input = 20'b00000010101011000110; // y = 0.1670854271356783 
#15 y_input = 20'b00000010110100110111; // y = 0.17663316582914557 
#15 y_input = 20'b00000010111110101001; // y = 0.18618090452261304 
#15 y_input = 20'b00000011001000011011; // y = 0.1957286432160803 
#15 y_input = 20'b00000011010010001100; // y = 0.20527638190954756 
#15 y_input = 20'b00000011011011111110; // y = 0.21482412060301503 
#15 y_input = 20'b00000011100101110000; // y = 0.2243718592964823 
#15 y_input = 20'b00000011101111100010; // y = 0.23391959798994977 
#15 y_input = 20'b00000011111001010011; // y = 0.24346733668341702 
#15 y_input = 20'b00000100000011000101; // y = 0.2530150753768843 
#15 y_input = 20'b00000100001100110111; // y = 0.26256281407035176 
#15 y_input = 20'b00000100010110101001; // y = 0.272110552763819 
#15 y_input = 20'b00000100100000011010; // y = 0.28165829145728627 
#15 y_input = 20'b00000100101010001100; // y = 0.29120603015075375 
#15 y_input = 20'b00000100110011111110; // y = 0.300753768844221 
#15 y_input = 20'b00000100111101101111; // y = 0.31030150753768826 
#15 y_input = 20'b00000101000111100001; // y = 0.31984924623115574 
#15 y_input = 20'b00000101010001010011; // y = 0.329396984924623 
#15 y_input = 20'b00000101011011000101; // y = 0.33894472361809047 
#15 y_input = 20'b00000101100100110110; // y = 0.3484924623115577 
#15 y_input = 20'b00000101101110101000; // y = 0.358040201005025 
#15 y_input = 20'b00000101111000011010; // y = 0.36758793969849246 
#15 y_input = 20'b00000110000010001011; // y = 0.3771356783919597 
#15 y_input = 20'b00000110001011111101; // y = 0.386683417085427 
#15 y_input = 20'b00000110010101101111; // y = 0.39623115577889445 
#15 y_input = 20'b00000110011111100001; // y = 0.4057788944723617 
#15 y_input = 20'b00000110101001010010; // y = 0.41532663316582896 
#15 y_input = 20'b00000110110011000100; // y = 0.42487437185929644 
#15 y_input = 20'b00000110111100110110; // y = 0.4344221105527637 
#15 y_input = 20'b00000111000110101000; // y = 0.44396984924623095 
#15 y_input = 20'b00000111010000011001; // y = 0.45351758793969843 
#15 y_input = 20'b00000111011010001011; // y = 0.4630653266331657 
#15 y_input = 20'b00000111100011111101; // y = 0.47261306532663316 
#15 y_input = 20'b00000111101101101110; // y = 0.4821608040201004 
#15 y_input = 20'b00000111110111100000; // y = 0.4917085427135677 
#15 y_input = 20'b00001000000001010010; // y = 0.5012562814070352 
#15 y_input = 20'b00001000001011000100; // y = 0.5108040201005024 
#15 y_input = 20'b00001000010100110101; // y = 0.5203517587939697 
#15 y_input = 20'b00001000011110100111; // y = 0.5298994974874371 
#15 y_input = 20'b00001000101000011001; // y = 0.5394472361809044 
#15 y_input = 20'b00001000110010001010; // y = 0.5489949748743717 
#15 y_input = 20'b00001000111011111100; // y = 0.5585427135678391 
#15 y_input = 20'b00001001000101101110; // y = 0.5680904522613064 
#15 y_input = 20'b00001001001111100000; // y = 0.5776381909547739 
#15 y_input = 20'b00001001011001010001; // y = 0.5871859296482411 
#15 y_input = 20'b00001001100011000011; // y = 0.5967336683417084 
#15 y_input = 20'b00001001101100110101; // y = 0.6062814070351759 
#15 y_input = 20'b00001001110110100110; // y = 0.6158291457286431 
#15 y_input = 20'b00001010000000011000; // y = 0.6253768844221104 
#15 y_input = 20'b00001010001010001010; // y = 0.6349246231155778 
#15 y_input = 20'b00001010010011111100; // y = 0.6444723618090451 
#15 y_input = 20'b00001010011101101101; // y = 0.6540201005025124 
#15 y_input = 20'b00001010100111011111; // y = 0.6635678391959798 
#15 y_input = 20'b00001010110001010001; // y = 0.6731155778894471 
#15 y_input = 20'b00001010111011000011; // y = 0.6826633165829143 
#15 y_input = 20'b00001011000100110100; // y = 0.6922110552763818 
#15 y_input = 20'b00001011001110100110; // y = 0.7017587939698491 
#15 y_input = 20'b00001011011000011000; // y = 0.7113065326633166 
#15 y_input = 20'b00001011100010001001; // y = 0.7208542713567838 
#15 y_input = 20'b00001011101011111011; // y = 0.7304020100502511 
#15 y_input = 20'b00001011110101101101; // y = 0.7399497487437185 
#15 y_input = 20'b00001011111111011111; // y = 0.7494974874371858 
#15 y_input = 20'b00001100001001010000; // y = 0.7590452261306531 
#15 y_input = 20'b00001100010011000010; // y = 0.7685929648241205 
#15 y_input = 20'b00001100011100110100; // y = 0.7781407035175878 
#15 y_input = 20'b00001100100110100101; // y = 0.787688442211055 
#15 y_input = 20'b00001100110000010111; // y = 0.7972361809045225 
#15 y_input = 20'b00001100111010001001; // y = 0.8067839195979898 
#15 y_input = 20'b00001101000011111011; // y = 0.816331658291457 
#15 y_input = 20'b00001101001101101100; // y = 0.8258793969849245 
#15 y_input = 20'b00001101010111011110; // y = 0.8354271356783918 
#15 y_input = 20'b00001101100001010000; // y = 0.8449748743718593 
#15 y_input = 20'b00001101101011000001; // y = 0.8545226130653265 
#15 y_input = 20'b00001101110100110011; // y = 0.8640703517587938 
#15 y_input = 20'b00001101111110100101; // y = 0.8736180904522612 
#15 y_input = 20'b00001110001000010111; // y = 0.8831658291457285 
#15 y_input = 20'b00001110010010001000; // y = 0.8927135678391958 
#15 y_input = 20'b00001110011011111010; // y = 0.9022613065326632 
#15 y_input = 20'b00001110100101101100; // y = 0.9118090452261305 
#15 y_input = 20'b00001110101111011110; // y = 0.9213567839195977 
#15 y_input = 20'b00001110111001001111; // y = 0.9309045226130652 
#15 y_input = 20'b00001111000011000001; // y = 0.9404522613065325 
#15 y_input = 20'b00001111001100110011; // y = 0.95 

      #15 $finish;
     end
endmodule
