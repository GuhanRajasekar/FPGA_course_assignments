`timescale 1ns / 1ps

module cordic_tanh_tb;
  reg  signed  [31:0] target_angle;
  reg clk,rst;
  wire signed [31:0] x_res;
  wire signed [31:0] y_res;
  wire signed [31:0] tanh_res;
  
  cordic_tanh w(.clk(clk),.rst(rst),.target_angle(target_angle), .x_res(x_res) , .y_res(y_res),.tanh_res(tanh_res));
  
  integer fh_tanh; // Variable for file handle
  
  always #2 clk = ~clk;
  
  /*
     for target angle the precision is 16 bits for integer part and 16 bits for the fractional part(Based on the look up table used)
     For the results, the precision is 16 bits for integer part and 16 bits for the fractional part
  */
  initial 
     begin
      #0 clk = 1'b0; rst = 1'b0; 
      #1 rst = 1'b1;
      fh_tanh = $fopen("F:/PhD_IISc/Coursework/Jan_2024/FPGA/FPGA_course_assignments/Mini_Project/Source_Code/Data/tanh_data.txt","w");
      $fmonitor(fh_tanh,"%b %d",tanh_res,target_angle);
      
//      #5 target_angle = 32'b00000000000000001000100011110101; // 0.535
//      #5 target_angle = 32'b11111111111111110111011100001011; // -0.535 (2's complement of 0.535)
//      #5 target_angle = {{14{1'b0}},2'b10,{16{1'b0}}}; // 2
//      #5 target_angle = {{16{1'b0}},16'b1100110011001100}; //0.8
//#15 target_angle = 32'b11111111111111110000000000000000; //-1.0 radians
#15 target_angle = 32'b11111111111111110000010100101100; //-0.9797979797979798 radians
#15 target_angle = 32'b11111111111111110000101001011000; //-0.9595959595959596 radians
#15 target_angle = 32'b11111111111111110000111110000100; //-0.9393939393939394 radians
#15 target_angle = 32'b11111111111111110001010010110000; //-0.9191919191919192 radians
#15 target_angle = 32'b11111111111111110001100111011100; //-0.898989898989899 radians
#15 target_angle = 32'b11111111111111110001111100001000; //-0.8787878787878788 radians
#15 target_angle = 32'b11111111111111110010010000110100; //-0.8585858585858586 radians
#15 target_angle = 32'b11111111111111110010100101100000; //-0.8383838383838383 radians
#15 target_angle = 32'b11111111111111110010111010001100; //-0.8181818181818181 radians
#15 target_angle = 32'b11111111111111110011001110111000; //-0.797979797979798 radians
#15 target_angle = 32'b11111111111111110011100011100100; //-0.7777777777777778 radians
#15 target_angle = 32'b11111111111111110011111000010000; //-0.7575757575757576 radians
#15 target_angle = 32'b11111111111111110100001100111100; //-0.7373737373737373 radians
#15 target_angle = 32'b11111111111111110100100001101000; //-0.7171717171717171 radians
#15 target_angle = 32'b11111111111111110100110110010100; //-0.696969696969697 radians
#15 target_angle = 32'b11111111111111110101001011000000; //-0.6767676767676767 radians
#15 target_angle = 32'b11111111111111110101011111101100; //-0.6565656565656566 radians
#15 target_angle = 32'b11111111111111110101110100011000; //-0.6363636363636364 radians
#15 target_angle = 32'b11111111111111110110001001000100; //-0.6161616161616161 radians
#15 target_angle = 32'b11111111111111110110011101110000; //-0.5959595959595959 radians
#15 target_angle = 32'b11111111111111110110110010011100; //-0.5757575757575757 radians
#15 target_angle = 32'b11111111111111110111000111001000; //-0.5555555555555556 radians
#15 target_angle = 32'b11111111111111110111011011110100; //-0.5353535353535352 radians
#15 target_angle = 32'b11111111111111110111110000100000; //-0.5151515151515151 radians
#15 target_angle = 32'b11111111111111111000000101001011; //-0.4949494949494949 radians
#15 target_angle = 32'b11111111111111111000011001110111; //-0.4747474747474747 radians
#15 target_angle = 32'b11111111111111111000101110100011; //-0.4545454545454545 radians
#15 target_angle = 32'b11111111111111111001000011001111; //-0.43434343434343425 radians
#15 target_angle = 32'b11111111111111111001010111111011; //-0.41414141414141414 radians
#15 target_angle = 32'b11111111111111111001101100100111; //-0.3939393939393939 radians
#15 target_angle = 32'b11111111111111111010000001010011; //-0.3737373737373737 radians
#15 target_angle = 32'b11111111111111111010010101111111; //-0.3535353535353535 radians
#15 target_angle = 32'b11111111111111111010101010101011; //-0.33333333333333326 radians
#15 target_angle = 32'b11111111111111111010111111010111; //-0.31313131313131304 radians
#15 target_angle = 32'b11111111111111111011010100000011; //-0.2929292929292928 radians
#15 target_angle = 32'b11111111111111111011101000101111; //-0.2727272727272727 radians
#15 target_angle = 32'b11111111111111111011111101011011; //-0.2525252525252525 radians
#15 target_angle = 32'b11111111111111111100010010000111; //-0.23232323232323226 radians
#15 target_angle = 32'b11111111111111111100100110110011; //-0.21212121212121204 radians
#15 target_angle = 32'b11111111111111111100111011011111; //-0.19191919191919182 radians
#15 target_angle = 32'b11111111111111111101010000001011; //-0.1717171717171716 radians
#15 target_angle = 32'b11111111111111111101100100110111; //-0.1515151515151515 radians
#15 target_angle = 32'b11111111111111111101111001100011; //-0.13131313131313127 radians
#15 target_angle = 32'b11111111111111111110001110001111; //-0.11111111111111105 radians
#15 target_angle = 32'b11111111111111111110100010111011; //-0.09090909090909083 radians
#15 target_angle = 32'b11111111111111111110110111100111; //-0.07070707070707061 radians
#15 target_angle = 32'b11111111111111111111001100010011; //-0.050505050505050386 radians
#15 target_angle = 32'b11111111111111111111100000111111; //-0.030303030303030276 radians
#15 target_angle = 32'b11111111111111111111110101101011; //-0.010101010101010055 radians
#15 target_angle = 32'b00000000000000000000001010010101; //0.010101010101010166 radians
#15 target_angle = 32'b00000000000000000000011111000001; //0.030303030303030498 radians
#15 target_angle = 32'b00000000000000000000110011101101; //0.05050505050505061 radians
#15 target_angle = 32'b00000000000000000001001000011001; //0.07070707070707072 radians
#15 target_angle = 32'b00000000000000000001011101000101; //0.09090909090909105 radians
#15 target_angle = 32'b00000000000000000001110001110001; //0.11111111111111116 radians
#15 target_angle = 32'b00000000000000000010000110011101; //0.1313131313131315 radians
#15 target_angle = 32'b00000000000000000010011011001001; //0.1515151515151516 radians
#15 target_angle = 32'b00000000000000000010101111110101; //0.1717171717171717 radians
#15 target_angle = 32'b00000000000000000011000100100001; //0.19191919191919204 radians
#15 target_angle = 32'b00000000000000000011011001001101; //0.21212121212121215 radians
#15 target_angle = 32'b00000000000000000011101101111001; //0.2323232323232325 radians
#15 target_angle = 32'b00000000000000000100000010100101; //0.2525252525252526 radians
#15 target_angle = 32'b00000000000000000100010111010001; //0.27272727272727293 radians
#15 target_angle = 32'b00000000000000000100101011111101; //0.29292929292929304 radians
#15 target_angle = 32'b00000000000000000101000000101001; //0.31313131313131315 radians
#15 target_angle = 32'b00000000000000000101010101010101; //0.3333333333333335 radians
#15 target_angle = 32'b00000000000000000101101010000001; //0.3535353535353536 radians
#15 target_angle = 32'b00000000000000000101111110101101; //0.3737373737373739 radians
#15 target_angle = 32'b00000000000000000110010011011001; //0.39393939393939403 radians
#15 target_angle = 32'b00000000000000000110101000000101; //0.41414141414141437 radians
#15 target_angle = 32'b00000000000000000110111100110001; //0.4343434343434345 radians
#15 target_angle = 32'b00000000000000000111010001011101; //0.4545454545454546 radians
#15 target_angle = 32'b00000000000000000111100110001001; //0.4747474747474749 radians
#15 target_angle = 32'b00000000000000000111111010110101; //0.49494949494949503 radians
#15 target_angle = 32'b00000000000000001000001111100000; //0.5151515151515154 radians
#15 target_angle = 32'b00000000000000001000100100001100; //0.5353535353535355 radians
#15 target_angle = 32'b00000000000000001000111000111000; //0.5555555555555556 radians
#15 target_angle = 32'b00000000000000001001001101100100; //0.5757575757575759 radians
#15 target_angle = 32'b00000000000000001001100010010000; //0.595959595959596 radians
#15 target_angle = 32'b00000000000000001001110110111100; //0.6161616161616164 radians
#15 target_angle = 32'b00000000000000001010001011101000; //0.6363636363636365 radians
#15 target_angle = 32'b00000000000000001010100000010100; //0.6565656565656568 radians
#15 target_angle = 32'b00000000000000001010110101000000; //0.6767676767676769 radians
#15 target_angle = 32'b00000000000000001011001001101100; //0.696969696969697 radians
#15 target_angle = 32'b00000000000000001011011110011000; //0.7171717171717173 radians
#15 target_angle = 32'b00000000000000001011110011000100; //0.7373737373737375 radians
#15 target_angle = 32'b00000000000000001100000111110000; //0.7575757575757578 radians
#15 target_angle = 32'b00000000000000001100011100011100; //0.7777777777777779 radians
#15 target_angle = 32'b00000000000000001100110001001000; //0.7979797979797982 radians
#15 target_angle = 32'b00000000000000001101000101110100; //0.8181818181818183 radians
#15 target_angle = 32'b00000000000000001101011010100000; //0.8383838383838385 radians
#15 target_angle = 32'b00000000000000001101101111001100; //0.8585858585858588 radians
#15 target_angle = 32'b00000000000000001110000011111000; //0.8787878787878789 radians
#15 target_angle = 32'b00000000000000001110011000100100; //0.8989898989898992 radians
#15 target_angle = 32'b00000000000000001110101101010000; //0.9191919191919193 radians
#15 target_angle = 32'b00000000000000001111000001111100; //0.9393939393939394 radians
#15 target_angle = 32'b00000000000000001111010110101000; //0.9595959595959598 radians
#15 target_angle = 32'b00000000000000001111101011010100; //0.9797979797979799 radians
#15 target_angle = 32'b00000000000000010000000000000000; //1.0 radians

$fclose(fh_tanh);

#15 $finish;
     end
endmodule
